//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      0416001 ���­� 0416225 ��¤�
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;

//Sign extended
always@(*) begin
	if(data_i[15]==1'b1) begin
		data_o[31:0] = {16'b1111111111111111 , data_i[15:0]};
	end
	else begin
		data_o[31:0] = {16'b0000000000000000 , data_i[15:0]};
	end
end          
endmodule      
     